module ac_tb;
	reg s1_tb, s2_tb, co2_tb, enable_tb;
	wire buzz_tb, led_tb;
	reg clk_tb;
	
	always #10;

	// always@(co2_tb)
	
endmodule
